module skullart (vccd1, vssd1);
 input vccd1;
 input vssd1;
endmodule
