magic
tech sky130A
timestamp 1670165111
<< metal1 >>
rect 4730 13300 6890 13570
rect 4460 13030 6890 13300
rect 3920 12490 7430 13030
rect 3650 11410 7700 12490
rect 3650 11140 4460 11410
rect 3650 10870 4190 11140
rect 3920 10600 4190 10870
rect 5270 10600 6080 11410
rect 6890 11140 7700 11410
rect 7160 10870 7700 11140
rect 7160 10600 7430 10870
rect 3920 10330 4460 10600
rect 5000 10330 6350 10600
rect 6890 10330 7430 10600
rect 3920 10060 5540 10330
rect 5810 10060 7160 10330
rect 4460 9790 5270 10060
rect 6080 9790 7160 10060
rect 4730 9250 6620 9790
rect 3110 8980 3920 9250
rect 4730 8980 5000 9250
rect 5270 8980 5540 9250
rect 5810 8980 6080 9250
rect 6350 8980 6620 9250
rect 7430 8980 8240 9250
rect 2840 8440 4190 8980
rect 7160 8440 8510 8980
rect 3110 8170 4730 8440
rect 6620 8170 8240 8440
rect 3920 7900 5000 8170
rect 6350 7900 7430 8170
rect 4460 7630 5540 7900
rect 5810 7630 6890 7900
rect 5000 7090 6350 7630
rect 4460 6820 5540 7090
rect 5810 6820 6890 7090
rect 3110 6550 5000 6820
rect 6350 6550 8510 6820
rect 2840 6280 4460 6550
rect 6890 6280 8510 6550
rect 2840 6010 3920 6280
rect 7430 6010 8510 6280
rect 2840 5740 3650 6010
rect 7700 5740 8510 6010
rect 3110 5470 3380 5740
rect 4730 5470 5000 5740
rect 5270 5470 5540 5740
rect 5810 5470 6080 5740
rect 6350 5470 6620 5740
rect 7970 5470 8240 5740
rect 4730 4930 6620 5470
rect 4460 4660 5270 4930
rect 6080 4660 7160 4930
rect 3920 4390 5540 4660
rect 5810 4390 7160 4660
rect 3920 4120 4460 4390
rect 5000 4120 6350 4390
rect 6890 4120 7430 4390
rect 3920 3850 4190 4120
rect 3650 3580 4190 3850
rect 3650 3310 4460 3580
rect 5270 3310 6080 4120
rect 7160 3850 7430 4120
rect 7160 3580 7700 3850
rect 6890 3310 7700 3580
rect 3650 2230 7700 3310
rect 3920 1690 7430 2230
rect 4460 1420 6890 1690
rect 4730 1150 6890 1420
<< metal4 >>
rect 1000 1000 1500 13570
rect 4730 13300 6890 13570
rect 4460 13030 6890 13300
rect 3920 12490 7430 13030
rect 3650 11410 7700 12490
rect 3650 11140 4460 11410
rect 3650 10870 4190 11140
rect 3920 10600 4190 10870
rect 5270 10600 6080 11410
rect 6890 11140 7700 11410
rect 7160 10870 7700 11140
rect 7160 10600 7430 10870
rect 3920 10330 4460 10600
rect 5000 10330 6350 10600
rect 6890 10330 7430 10600
rect 3920 10060 5540 10330
rect 5810 10060 7160 10330
rect 4460 9790 5270 10060
rect 6080 9790 7160 10060
rect 4730 9250 6620 9790
rect 3110 8980 3920 9250
rect 4730 8980 5000 9250
rect 5270 8980 5540 9250
rect 5810 8980 6080 9250
rect 6350 8980 6620 9250
rect 7430 8980 8240 9250
rect 2840 8440 4190 8980
rect 7160 8440 8510 8980
rect 3110 8170 4730 8440
rect 6620 8170 8240 8440
rect 3920 7900 5000 8170
rect 6350 7900 7430 8170
rect 4460 7630 5540 7900
rect 5810 7630 6890 7900
rect 5000 7090 6350 7630
rect 4460 6820 5540 7090
rect 5810 6820 6890 7090
rect 3110 6550 5000 6820
rect 6350 6550 8510 6820
rect 2840 6280 4460 6550
rect 6890 6280 8510 6550
rect 2840 6010 3920 6280
rect 7430 6010 8510 6280
rect 2840 5740 3650 6010
rect 7700 5740 8510 6010
rect 3110 5470 3380 5740
rect 4730 5470 5000 5740
rect 5270 5470 5540 5740
rect 5810 5470 6080 5740
rect 6350 5470 6620 5740
rect 7970 5470 8240 5740
rect 4730 4930 6620 5470
rect 4460 4660 5270 4930
rect 6080 4660 7160 4930
rect 3920 4390 5540 4660
rect 5810 4390 7160 4660
rect 3920 4120 4460 4390
rect 5000 4120 6350 4390
rect 6890 4120 7430 4390
rect 3920 3850 4190 4120
rect 3650 3580 4190 3850
rect 3650 3310 4460 3580
rect 5270 3310 6080 4120
rect 7160 3850 7430 4120
rect 7160 3580 7700 3850
rect 6890 3310 7700 3580
rect 3650 2230 7700 3310
rect 3920 1690 7430 2230
rect 4460 1420 6890 1690
rect 4730 1150 6890 1420
rect 9500 1000 10000 13570
<< labels >>
flabel metal4 s 9500 6500 10000 7500 0 FreeSans 240 0 0 0 vssd1
port 1 nsew ground bidirectional abutment
flabel metal4 s 1000 6500 1500 7500 0 FreeSans 240 0 0 0 vccd1
port 2 nsew power bidirectional abutment
<< end >>
