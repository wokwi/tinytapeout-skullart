magic
tech sky130A
timestamp 1670241224
<< metal1 >>
rect 7030 16150 9190 16420
rect 6760 15880 9190 16150
rect 6220 15340 9730 15880
rect 5950 14260 10000 15340
rect 5950 13990 6760 14260
rect 5950 13720 6490 13990
rect 6220 13450 6490 13720
rect 7570 13450 8380 14260
rect 9190 13990 10000 14260
rect 9460 13720 10000 13990
rect 9460 13450 9730 13720
rect 6220 13180 6760 13450
rect 7300 13180 8650 13450
rect 9190 13180 9730 13450
rect 6220 12910 7840 13180
rect 8110 12910 9460 13180
rect 6760 12640 7570 12910
rect 8380 12640 9460 12910
rect 7030 12100 8920 12640
rect 5410 11830 6220 12100
rect 7030 11830 7300 12100
rect 7570 11830 7840 12100
rect 8110 11830 8380 12100
rect 8650 11830 8920 12100
rect 9730 11830 10540 12100
rect 5140 11290 6490 11830
rect 9460 11290 10810 11830
rect 5410 11020 7030 11290
rect 8920 11020 10540 11290
rect 6220 10750 7300 11020
rect 8650 10750 9730 11020
rect 6760 10480 7840 10750
rect 8110 10480 9190 10750
rect 7300 9940 8650 10480
rect 6760 9670 7840 9940
rect 8110 9670 9190 9940
rect 5410 9400 7300 9670
rect 8650 9400 10810 9670
rect 5140 9130 6760 9400
rect 9190 9130 10810 9400
rect 5140 8860 6220 9130
rect 9730 8860 10810 9130
rect 5140 8590 5950 8860
rect 10000 8590 10810 8860
rect 5410 8320 5680 8590
rect 7030 8320 7300 8590
rect 7570 8320 7840 8590
rect 8110 8320 8380 8590
rect 8650 8320 8920 8590
rect 10270 8320 10540 8590
rect 7030 7780 8920 8320
rect 6760 7510 7570 7780
rect 8380 7510 9460 7780
rect 6220 7240 7840 7510
rect 8110 7240 9460 7510
rect 6220 6970 6760 7240
rect 7300 6970 8650 7240
rect 9190 6970 9730 7240
rect 6220 6700 6490 6970
rect 5950 6430 6490 6700
rect 5950 6160 6760 6430
rect 7570 6160 8380 6970
rect 9460 6700 9730 6970
rect 9460 6430 10000 6700
rect 9190 6160 10000 6430
rect 5950 5080 10000 6160
rect 6220 4540 9730 5080
rect 6760 4270 9190 4540
rect 7030 4000 9190 4270
rect 3400 3100 4200 3200
rect 4700 3100 4800 3200
rect 3300 3000 4200 3100
rect 4600 3000 4800 3100
rect 3200 2400 3500 3000
rect 3900 2800 4200 3000
rect 3900 2700 4100 2800
rect 3900 2600 4000 2700
rect 4500 2600 4800 3000
rect 5200 3100 5300 3200
rect 5100 3000 5400 3100
rect 5000 2900 5400 3000
rect 4900 2800 5300 2900
rect 4900 2700 5200 2800
rect 4900 2600 5100 2700
rect 4500 2500 5100 2600
rect 4400 2400 5000 2500
rect 3000 2300 4200 2400
rect 4300 2300 5000 2400
rect 3100 2200 4200 2300
rect 3400 1900 3500 2000
rect 3300 1800 3500 1900
rect 3900 1800 4200 2200
rect 4500 2200 5100 2300
rect 3200 1700 4100 1800
rect 3100 1600 4000 1700
rect 4500 1600 4800 2200
rect 4900 2100 5100 2200
rect 4900 2000 5200 2100
rect 4900 1900 5300 2000
rect 5000 1800 5400 1900
rect 5100 1700 5400 1800
rect 5500 1800 5800 3200
rect 6200 3100 6300 3200
rect 6800 3100 6900 3200
rect 7800 3100 7900 3200
rect 9000 3100 9800 3200
rect 10300 3100 11100 3200
rect 6200 3000 6400 3100
rect 6700 3000 6900 3100
rect 7700 3000 7900 3100
rect 8900 3000 9800 3100
rect 10200 3000 11100 3100
rect 11600 3000 11900 3200
rect 6200 1800 6500 3000
rect 6600 1800 6900 3000
rect 7400 1800 7500 1900
rect 5500 1700 6400 1800
rect 6600 1700 7100 1800
rect 7300 1700 7500 1800
rect 5200 1600 5300 1700
rect 5500 1600 6300 1700
rect 6600 1600 7500 1700
rect 7600 1800 7900 3000
rect 8800 2500 9100 3000
rect 9500 2800 9800 3000
rect 9500 2700 9700 2800
rect 9500 2600 9600 2700
rect 10100 2500 10400 3000
rect 10800 2800 11100 3000
rect 11200 2900 12200 3000
rect 11300 2800 12300 2900
rect 10800 2700 11000 2800
rect 11500 2700 12300 2800
rect 10800 2600 10900 2700
rect 8700 2400 9400 2500
rect 10000 2400 10700 2500
rect 8600 2300 9400 2400
rect 9900 2300 10700 2400
rect 8400 1800 8500 1900
rect 7600 1700 8100 1800
rect 8300 1700 8500 1800
rect 7600 1600 8500 1700
rect 8800 1600 9100 2300
rect 10100 1800 10400 2300
rect 10800 2100 10900 2200
rect 10800 2000 11000 2100
rect 10800 1800 11100 2000
rect 10100 1600 11100 1800
rect 11600 1800 11900 2700
rect 12100 2600 12300 2700
rect 12200 2500 12300 2600
rect 11600 1700 12100 1800
rect 11500 1600 12000 1700
rect 4500 1500 4600 1600
rect 6600 1500 6700 1600
rect 7600 1500 7700 1600
<< obsm2 >>
rect 5000 4000 11000 17000
rect 2500 1000 13000 4000
<< obsm3 >>
rect 5000 4000 11000 17000
rect 2500 1000 13000 4000
<< metal4 >>
rect 1000 1000 1500 17000
rect 7030 16150 9190 16420
rect 6760 15880 9190 16150
rect 6220 15340 9730 15880
rect 5950 14260 10000 15340
rect 5950 13990 6760 14260
rect 5950 13720 6490 13990
rect 6220 13450 6490 13720
rect 7570 13450 8380 14260
rect 9190 13990 10000 14260
rect 9460 13720 10000 13990
rect 9460 13450 9730 13720
rect 6220 13180 6760 13450
rect 7300 13180 8650 13450
rect 9190 13180 9730 13450
rect 6220 12910 7840 13180
rect 8110 12910 9460 13180
rect 6760 12640 7570 12910
rect 8380 12640 9460 12910
rect 7030 12100 8920 12640
rect 5410 11830 6220 12100
rect 7030 11830 7300 12100
rect 7570 11830 7840 12100
rect 8110 11830 8380 12100
rect 8650 11830 8920 12100
rect 9730 11830 10540 12100
rect 5140 11290 6490 11830
rect 9460 11290 10810 11830
rect 5410 11020 7030 11290
rect 8920 11020 10540 11290
rect 6220 10750 7300 11020
rect 8650 10750 9730 11020
rect 6760 10480 7840 10750
rect 8110 10480 9190 10750
rect 7300 9940 8650 10480
rect 6760 9670 7840 9940
rect 8110 9670 9190 9940
rect 5410 9400 7300 9670
rect 8650 9400 10810 9670
rect 5140 9130 6760 9400
rect 9190 9130 10810 9400
rect 5140 8860 6220 9130
rect 9730 8860 10810 9130
rect 5140 8590 5950 8860
rect 10000 8590 10810 8860
rect 5410 8320 5680 8590
rect 7030 8320 7300 8590
rect 7570 8320 7840 8590
rect 8110 8320 8380 8590
rect 8650 8320 8920 8590
rect 10270 8320 10540 8590
rect 7030 7780 8920 8320
rect 6760 7510 7570 7780
rect 8380 7510 9460 7780
rect 6220 7240 7840 7510
rect 8110 7240 9460 7510
rect 6220 6970 6760 7240
rect 7300 6970 8650 7240
rect 9190 6970 9730 7240
rect 6220 6700 6490 6970
rect 5950 6430 6490 6700
rect 5950 6160 6760 6430
rect 7570 6160 8380 6970
rect 9460 6700 9730 6970
rect 9460 6430 10000 6700
rect 9190 6160 10000 6430
rect 5950 5080 10000 6160
rect 6220 4540 9730 5080
rect 6760 4270 9190 4540
rect 7030 4000 9190 4270
rect 3400 3100 4200 3200
rect 4700 3100 4800 3200
rect 3300 3000 4200 3100
rect 4600 3000 4800 3100
rect 3200 2400 3500 3000
rect 3900 2800 4200 3000
rect 3900 2700 4100 2800
rect 3900 2600 4000 2700
rect 4500 2600 4800 3000
rect 5200 3100 5300 3200
rect 5100 3000 5400 3100
rect 5000 2900 5400 3000
rect 4900 2800 5300 2900
rect 4900 2700 5200 2800
rect 4900 2600 5100 2700
rect 4500 2500 5100 2600
rect 4400 2400 5000 2500
rect 3000 2300 4200 2400
rect 4300 2300 5000 2400
rect 3100 2200 4200 2300
rect 3400 1900 3500 2000
rect 3300 1800 3500 1900
rect 3900 1800 4200 2200
rect 4500 2200 5100 2300
rect 3200 1700 4100 1800
rect 3100 1600 4000 1700
rect 4500 1600 4800 2200
rect 4900 2100 5100 2200
rect 4900 2000 5200 2100
rect 4900 1900 5300 2000
rect 5000 1800 5400 1900
rect 5100 1700 5400 1800
rect 5500 1800 5800 3200
rect 6200 3100 6300 3200
rect 6800 3100 6900 3200
rect 7800 3100 7900 3200
rect 9000 3100 9800 3200
rect 10300 3100 11100 3200
rect 6200 3000 6400 3100
rect 6700 3000 6900 3100
rect 7700 3000 7900 3100
rect 8900 3000 9800 3100
rect 10200 3000 11100 3100
rect 11600 3000 11900 3200
rect 6200 1800 6500 3000
rect 6600 1800 6900 3000
rect 7400 1800 7500 1900
rect 5500 1700 6400 1800
rect 6600 1700 7100 1800
rect 7300 1700 7500 1800
rect 5200 1600 5300 1700
rect 5500 1600 6300 1700
rect 6600 1600 7500 1700
rect 7600 1800 7900 3000
rect 8800 2500 9100 3000
rect 9500 2800 9800 3000
rect 9500 2700 9700 2800
rect 9500 2600 9600 2700
rect 10100 2500 10400 3000
rect 10800 2800 11100 3000
rect 11200 2900 12200 3000
rect 11300 2800 12300 2900
rect 10800 2700 11000 2800
rect 11500 2700 12300 2800
rect 10800 2600 10900 2700
rect 8700 2400 9400 2500
rect 10000 2400 10700 2500
rect 8600 2300 9400 2400
rect 9900 2300 10700 2400
rect 8400 1800 8500 1900
rect 7600 1700 8100 1800
rect 8300 1700 8500 1800
rect 7600 1600 8500 1700
rect 8800 1600 9100 2300
rect 10100 1800 10400 2300
rect 10800 2100 10900 2200
rect 10800 2000 11000 2100
rect 10800 1800 11100 2000
rect 10100 1600 11100 1800
rect 11600 1800 11900 2700
rect 12100 2600 12300 2700
rect 12200 2500 12300 2600
rect 11600 1700 12100 1800
rect 11500 1600 12000 1700
rect 4500 1500 4600 1600
rect 6600 1500 6700 1600
rect 7600 1500 7700 1600
rect 14500 1000 15000 17000
<< labels >>
flabel metal4 s 14500 16500 15000 17000 0 FreeSans 240 0 0 0 vssd1
port 1 nsew ground bidirectional abutment
flabel metal4 s 1000 16500 1500 17000 0 FreeSans 240 0 0 0 vccd1
port 2 nsew power bidirectional abutment
<< end >>
