magic
tech sky130A
timestamp 1670235840
<< metal1 >>
rect 7030 14950 9190 15220
rect 6760 14680 9190 14950
rect 6220 14140 9730 14680
rect 5950 13060 10000 14140
rect 5950 12790 6760 13060
rect 5950 12520 6490 12790
rect 6220 12250 6490 12520
rect 7570 12250 8380 13060
rect 9190 12790 10000 13060
rect 9460 12520 10000 12790
rect 9460 12250 9730 12520
rect 6220 11980 6760 12250
rect 7300 11980 8650 12250
rect 9190 11980 9730 12250
rect 6220 11710 7840 11980
rect 8110 11710 9460 11980
rect 6760 11440 7570 11710
rect 8380 11440 9460 11710
rect 7030 10900 8920 11440
rect 5410 10630 6220 10900
rect 7030 10630 7300 10900
rect 7570 10630 7840 10900
rect 8110 10630 8380 10900
rect 8650 10630 8920 10900
rect 9730 10630 10540 10900
rect 5140 10090 6490 10630
rect 9460 10090 10810 10630
rect 5410 9820 7030 10090
rect 8920 9820 10540 10090
rect 6220 9550 7300 9820
rect 8650 9550 9730 9820
rect 6760 9280 7840 9550
rect 8110 9280 9190 9550
rect 7300 8740 8650 9280
rect 6760 8470 7840 8740
rect 8110 8470 9190 8740
rect 5410 8200 7300 8470
rect 8650 8200 10810 8470
rect 5140 7930 6760 8200
rect 9190 7930 10810 8200
rect 5140 7660 6220 7930
rect 9730 7660 10810 7930
rect 5140 7390 5950 7660
rect 10000 7390 10810 7660
rect 5410 7120 5680 7390
rect 7030 7120 7300 7390
rect 7570 7120 7840 7390
rect 8110 7120 8380 7390
rect 8650 7120 8920 7390
rect 10270 7120 10540 7390
rect 7030 6580 8920 7120
rect 6760 6310 7570 6580
rect 8380 6310 9460 6580
rect 6220 6040 7840 6310
rect 8110 6040 9460 6310
rect 6220 5770 6760 6040
rect 7300 5770 8650 6040
rect 9190 5770 9730 6040
rect 6220 5500 6490 5770
rect 5950 5230 6490 5500
rect 5950 4960 6760 5230
rect 7570 4960 8380 5770
rect 9460 5500 9730 5770
rect 9460 5230 10000 5500
rect 9190 4960 10000 5230
rect 5950 3880 10000 4960
rect 6220 3340 9730 3880
rect 6760 3070 9190 3340
rect 7030 2800 9190 3070
<< metal4 >>
rect 1000 1000 1500 17000
rect 7030 14950 9190 15220
rect 6760 14680 9190 14950
rect 6220 14140 9730 14680
rect 5950 13060 10000 14140
rect 5950 12790 6760 13060
rect 5950 12520 6490 12790
rect 6220 12250 6490 12520
rect 7570 12250 8380 13060
rect 9190 12790 10000 13060
rect 9460 12520 10000 12790
rect 9460 12250 9730 12520
rect 6220 11980 6760 12250
rect 7300 11980 8650 12250
rect 9190 11980 9730 12250
rect 6220 11710 7840 11980
rect 8110 11710 9460 11980
rect 6760 11440 7570 11710
rect 8380 11440 9460 11710
rect 7030 10900 8920 11440
rect 5410 10630 6220 10900
rect 7030 10630 7300 10900
rect 7570 10630 7840 10900
rect 8110 10630 8380 10900
rect 8650 10630 8920 10900
rect 9730 10630 10540 10900
rect 5140 10090 6490 10630
rect 9460 10090 10810 10630
rect 5410 9820 7030 10090
rect 8920 9820 10540 10090
rect 6220 9550 7300 9820
rect 8650 9550 9730 9820
rect 6760 9280 7840 9550
rect 8110 9280 9190 9550
rect 7300 8740 8650 9280
rect 6760 8470 7840 8740
rect 8110 8470 9190 8740
rect 5410 8200 7300 8470
rect 8650 8200 10810 8470
rect 5140 7930 6760 8200
rect 9190 7930 10810 8200
rect 5140 7660 6220 7930
rect 9730 7660 10810 7930
rect 5140 7390 5950 7660
rect 10000 7390 10810 7660
rect 5410 7120 5680 7390
rect 7030 7120 7300 7390
rect 7570 7120 7840 7390
rect 8110 7120 8380 7390
rect 8650 7120 8920 7390
rect 10270 7120 10540 7390
rect 7030 6580 8920 7120
rect 6760 6310 7570 6580
rect 8380 6310 9460 6580
rect 6220 6040 7840 6310
rect 8110 6040 9460 6310
rect 6220 5770 6760 6040
rect 7300 5770 8650 6040
rect 9190 5770 9730 6040
rect 6220 5500 6490 5770
rect 5950 5230 6490 5500
rect 5950 4960 6760 5230
rect 7570 4960 8380 5770
rect 9460 5500 9730 5770
rect 9460 5230 10000 5500
rect 9190 4960 10000 5230
rect 5950 3880 10000 4960
rect 6220 3340 9730 3880
rect 6760 3070 9190 3340
rect 7030 2800 9190 3070
rect 14500 1000 15000 17000
<< obsm2 >>
rect 5000 2500 11000 15500
<< obsm3 >>
rect 5000 2500 11000 15500
<< labels >>
flabel metal4 s 14500 16500 15000 17000 0 FreeSans 240 0 0 0 vssd1
port 1 nsew ground bidirectional abutment
flabel metal4 s 1000 16500 1500 17000 0 FreeSans 240 0 0 0 vccd1
port 2 nsew power bidirectional abutment
<< end >>
