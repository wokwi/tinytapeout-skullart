`default_nettype none

module skullart(
);
endmodule
